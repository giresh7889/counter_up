resh very good boy
